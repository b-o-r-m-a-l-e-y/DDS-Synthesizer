module sin_lut(clk, addr, q);
input clk;
input addr


endmodule